-------------------------------------------------------------------------------
-- COPYRIGHT (c) SOLECTRIX GmbH, Germany, 2017            All rights reserved
--
-- The copyright to the document(s) herein is the property of SOLECTRIX GmbH
-- The document(s) may be used AND/OR copied only with the written permission
-- from SOLECTRIX GmbH or in accordance with the terms/conditions stipulated
-- in the agreement/contract under which the document(s) have been supplied
-------------------------------------------------------------------------------
--*
--* @short INTERCON
--*        Generated by TCL script gen_intercon.tcl. Do not edit this file.
--* @author wrupprecht
--*
-------------------------------------------------------------------------------
-- for defines see wbi_test.sxl
--
-- Generated Tue Jun 20 15:35:45 CEST 2017
--
-- Wishbone masters:
--   wbm_1
--   wbm_2
--
-- Wishbone slaves:
--   wbs_1
--     baseaddr 0x00000000 - size 0x00000100
--   wbs_2
--     baseaddr 0x00000200 - size 0x00000010
--   wbs_3
--     baseaddr 0x00100000 - size 0x00001000
--
-- Intercon type: SharedBus
--
-------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

LIBRARY rtl_lib;

ENTITY wbi_test IS
  PORT (
    -- wishbone master port(s)
    -- wbm_1
    i_wbm_1_o_cyc       : IN  STD_LOGIC;
    i_wbm_1_o_stb       : IN  STD_LOGIC;
    i_wbm_1_o_we        : IN  STD_LOGIC;
    i_wbm_1_o_sel       : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    i_wbm_1_o_addr      : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
    i_wbm_1_o_data      : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
    o_wbm_1_i_data      : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    o_wbm_1_i_ack       : OUT STD_LOGIC;
    o_wbm_1_i_rty       : OUT STD_LOGIC;
    o_wbm_1_i_err       : OUT STD_LOGIC;
    -- wbm_2
    i_wbm_2_o_cyc       : IN  STD_LOGIC;
    i_wbm_2_o_stb       : IN  STD_LOGIC;
    i_wbm_2_o_we        : IN  STD_LOGIC;
    i_wbm_2_o_sel       : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    i_wbm_2_o_addr      : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
    i_wbm_2_o_data      : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
    o_wbm_2_i_data      : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    o_wbm_2_i_ack       : OUT STD_LOGIC;
    o_wbm_2_i_rty       : OUT STD_LOGIC;
    o_wbm_2_i_err       : OUT STD_LOGIC;
    -- wishbone slave port(s)
    -- wbs_1
    o_wbs_1_i_cyc       : OUT STD_LOGIC;
    o_wbs_1_i_stb       : OUT STD_LOGIC;
    o_wbs_1_i_we        : OUT STD_LOGIC;
    o_wbs_1_i_sel       : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    o_wbs_1_i_addr      : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    o_wbs_1_i_data      : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    i_wbs_1_o_data      : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
    i_wbs_1_o_ack       : IN  STD_LOGIC;
    i_wbs_1_o_rty       : IN  STD_LOGIC;
    i_wbs_1_o_err       : IN  STD_LOGIC;
    -- wbs_2
    o_wbs_2_i_cyc       : OUT STD_LOGIC;
    o_wbs_2_i_stb       : OUT STD_LOGIC;
    o_wbs_2_i_sel       : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    o_wbs_2_i_addr      : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    i_wbs_2_o_data      : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
    i_wbs_2_o_ack       : IN  STD_LOGIC;
    i_wbs_2_o_rty       : IN  STD_LOGIC;
    i_wbs_2_o_err       : IN  STD_LOGIC;
    -- wbs_3
    o_wbs_3_i_cyc       : OUT STD_LOGIC;
    o_wbs_3_i_stb       : OUT STD_LOGIC;
    o_wbs_3_i_we        : OUT STD_LOGIC;
    o_wbs_3_i_sel       : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    o_wbs_3_i_addr      : OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
    o_wbs_3_i_data      : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    i_wbs_3_o_data      : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
    i_wbs_3_o_ack       : IN  STD_LOGIC;
    i_wbs_3_o_rty       : IN  STD_LOGIC;
    i_wbs_3_o_err       : IN  STD_LOGIC;
    -- clock and reset
    clk                 : IN  STD_LOGIC;
    rst_n               : IN  STD_LOGIC := '1');
END ENTITY wbi_test;

-------------------------------------------------------------------------------

ARCHITECTURE rtl OF wbi_test IS

  FUNCTION "AND" (
    le : STD_LOGIC_VECTOR;
    ri : STD_LOGIC)
    RETURN STD_LOGIC_VECTOR IS
    VARIABLE v_result : STD_LOGIC_VECTOR(le'RANGE);
  BEGIN
    FOR i IN le'RANGE LOOP
      v_result(i) := le(i) AND ri;
    END LOOP;
    RETURN v_result;
  END FUNCTION "AND";

  SIGNAL s_wbm_1_bg        : STD_LOGIC; -- bus grant
  SIGNAL s_wbm_2_bg        : STD_LOGIC; -- bus grant
  SIGNAL s_wbs_1_ss        : STD_LOGIC; -- slave select
  SIGNAL s_wbs_2_ss        : STD_LOGIC; -- slave select
  SIGNAL s_wbs_3_ss        : STD_LOGIC; -- slave select

BEGIN  -- rtl

  arbiter_sharedbus : BLOCK
    SIGNAL s_wbm_1_bg_1      : STD_LOGIC;
    SIGNAL s_wbm_1_bb_1      : STD_LOGIC;
    SIGNAL s_wbm_1_bg_2      : STD_LOGIC;
    SIGNAL s_wbm_1_bb_2      : STD_LOGIC;
    SIGNAL s_wbm_1_bg_q      : STD_LOGIC;
    SIGNAL s_wbm_2_bg_1      : STD_LOGIC;
    SIGNAL s_wbm_2_bb_1      : STD_LOGIC;
    SIGNAL s_wbm_2_bg_2      : STD_LOGIC;
    SIGNAL s_wbm_2_bb_2      : STD_LOGIC;
    SIGNAL s_wbm_2_bg_q      : STD_LOGIC;
    SIGNAL s_wbm_1_traffic_ctrl_limit : STD_LOGIC;
    SIGNAL s_wbm_2_traffic_ctrl_limit : STD_LOGIC;
    SIGNAL s_ack             : STD_LOGIC;
    SIGNAL s_ce              : STD_LOGIC;
    SIGNAL s_idle            : STD_LOGIC;
  BEGIN -- arbiter
    s_ack <= i_wbs_1_o_ack OR i_wbs_2_o_ack OR i_wbs_3_o_ack;

    wb_traffic_supervision_1 : ENTITY rtl_lib.wb_traffic_supervision
      GENERIC MAP (
        g_priority     => 1,
        g_tot_priority => 2)
      PORT MAP (
        i_bg            => s_wbm_1_bg,
        i_ce            => s_ce,
        o_traffic_limit => s_wbm_1_traffic_ctrl_limit,
        clk             => clk,
        rst_n           => rst_n);

    wb_traffic_supervision_2 : ENTITY rtl_lib.wb_traffic_supervision
      GENERIC MAP (
        g_priority     => 1,
        g_tot_priority => 2)
      PORT MAP (
        i_bg            => s_wbm_2_bg,
        i_ce            => s_ce,
        o_traffic_limit => s_wbm_2_traffic_ctrl_limit,
        clk             => clk,
        rst_n           => rst_n);

    PROCESS (clk, rst_n)
    BEGIN
      IF (rst_n = '0') THEN
        s_wbm_1_bg_q <= '0';
      ELSIF (clk'EVENT AND clk = '1') THEN
        IF (s_wbm_1_bg_q = '0') THEN
          s_wbm_1_bg_q <= s_wbm_1_bg;
        ELSIF (s_ack = '1') THEN
          s_wbm_1_bg_q <= '0';
        ELSIF (i_wbm_1_o_cyc = '0') THEN
          s_wbm_1_bg_q <= '0';
        END IF;
      END IF;
    END PROCESS;

    PROCESS (clk, rst_n)
    BEGIN
      IF (rst_n = '0') THEN
        s_wbm_2_bg_q <= '0';
      ELSIF (clk'EVENT AND clk = '1') THEN
        IF (s_wbm_2_bg_q = '0') THEN
          s_wbm_2_bg_q <= s_wbm_2_bg;
        ELSIF (s_ack = '1') THEN
          s_wbm_2_bg_q <= '0';
        ELSIF (i_wbm_2_o_cyc = '0') THEN
          s_wbm_2_bg_q <= '0';
        END IF;
      END IF;
    END PROCESS;

    s_idle <= '1' WHEN (s_wbm_1_bg_q = '0' AND s_wbm_2_bg_q = '0') ELSE '0';
    s_wbm_1_bg_1 <= '1' WHEN (s_idle = '1' AND i_wbm_1_o_cyc = '1' AND s_wbm_1_traffic_ctrl_limit = '0') ELSE '0';
    s_wbm_1_bb_1 <= '1' WHEN (s_wbm_1_bg_1 = '1') ELSE '0';
    s_wbm_2_bg_1 <= '1' WHEN (s_idle = '1' AND i_wbm_2_o_cyc = '1' AND s_wbm_2_traffic_ctrl_limit = '0' AND s_wbm_1_bb_1 = '0') ELSE '0';
    s_wbm_2_bb_1 <= '1' WHEN (s_wbm_2_bg_1 = '1' OR s_wbm_1_bb_1 = '1') ELSE '0';
    s_wbm_1_bg_2 <= '1' WHEN (s_idle = '1' AND s_wbm_2_bb_1 = '0' AND i_wbm_1_o_cyc = '1') ELSE '0';
    s_wbm_1_bb_2 <= '1' WHEN (s_wbm_1_bg_2 = '1' OR s_wbm_2_bb_1 = '1') ELSE '0';
    s_wbm_2_bg_2 <= '1' WHEN (s_idle = '1' AND s_wbm_1_bb_2 = '0' AND i_wbm_2_o_cyc = '1') ELSE '0';
    s_wbm_2_bb_2 <= '1' WHEN (s_wbm_2_bg_2 = '1' OR s_wbm_1_bb_2 = '1') ELSE '0';
    s_wbm_1_bg   <= s_wbm_1_bg_q OR s_wbm_1_bg_1 OR s_wbm_1_bg_2;
    s_wbm_2_bg   <= s_wbm_2_bg_q OR s_wbm_2_bg_1 OR s_wbm_2_bg_2;
    s_ce <= i_wbm_1_o_cyc OR i_wbm_2_o_cyc WHEN (s_idle = '1') ELSE '0';
  END BLOCK arbiter_sharedbus;

  decoder : BLOCK
    SIGNAL s_addr : STD_LOGIC_VECTOR(31 DOWNTO 0);
  BEGIN
    s_addr <= (i_wbm_1_o_addr AND s_wbm_1_bg) OR (i_wbm_2_o_addr AND s_wbm_2_bg);
    s_wbs_1_ss <=
      '1' WHEN (s_addr(31 DOWNTO 8) = "000000000000000000000000") ELSE '0';
    s_wbs_2_ss <=
      '1' WHEN (s_addr(31 DOWNTO 4) = "0000000000000000000000100000") ELSE '0';
    s_wbs_3_ss <=
      '1' WHEN (s_addr(31 DOWNTO 12) = "00000000000100000000") ELSE '0';

    o_wbs_1_i_addr      <= s_addr(7 DOWNTO 0);
    o_wbs_2_i_addr      <= s_addr(3 DOWNTO 0);
    o_wbs_3_i_addr      <= s_addr(19 DOWNTO 0);
  END BLOCK decoder;

  mux : BLOCK
    SIGNAL s_cyc      : STD_LOGIC;
    SIGNAL s_stb      : STD_LOGIC;
    SIGNAL s_sel      : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL s_we       : STD_LOGIC;
    SIGNAL s_data_m2s : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL s_data_s2m : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL s_ack      : STD_LOGIC;
    SIGNAL s_rty      : STD_LOGIC;
    SIGNAL s_err      : STD_LOGIC;
  BEGIN
    -- cyc
    s_cyc <= (i_wbm_1_o_cyc AND s_wbm_1_bg) OR (i_wbm_2_o_cyc AND s_wbm_2_bg);
    o_wbs_1_i_cyc       <= s_cyc AND s_wbs_1_ss;
    o_wbs_2_i_cyc       <= s_cyc AND s_wbs_2_ss;
    o_wbs_3_i_cyc       <= s_cyc AND s_wbs_3_ss;
    -- stb
    s_stb <= (i_wbm_1_o_stb AND s_wbm_1_bg) OR (i_wbm_2_o_stb AND s_wbm_2_bg);
    o_wbs_1_i_stb       <= s_stb AND s_wbs_1_ss;
    o_wbs_2_i_stb       <= s_stb AND s_wbs_2_ss;
    o_wbs_3_i_stb       <= s_stb AND s_wbs_3_ss;
    -- sel
    s_sel <= (i_wbm_1_o_sel AND s_wbm_1_bg) OR (i_wbm_2_o_sel AND s_wbm_2_bg);
    o_wbs_1_i_sel       <= s_sel;
    o_wbs_2_i_sel       <= s_sel;
    o_wbs_3_i_sel       <= s_sel;
    -- we
    s_we <= (i_wbm_1_o_we AND s_wbm_1_bg) OR (i_wbm_2_o_we AND s_wbm_2_bg);
    o_wbs_1_i_we        <= s_we;
    o_wbs_3_i_we        <= s_we;
    -- data m2s
    s_data_m2s <= (i_wbm_1_o_data AND s_wbm_1_bg) OR (i_wbm_2_o_data AND s_wbm_2_bg);
    o_wbs_1_i_data      <= s_data_m2s;
    o_wbs_3_i_data      <= s_data_m2s;
    -- data s2m
    s_data_s2m <= (i_wbs_1_o_data AND s_wbs_1_ss) OR (i_wbs_2_o_data AND s_wbs_2_ss) OR (i_wbs_3_o_data AND s_wbs_3_ss);
    o_wbm_1_i_data      <= s_data_s2m;
    o_wbm_2_i_data      <= s_data_s2m;
    -- ack
    s_ack <= i_wbs_1_o_ack OR i_wbs_2_o_ack OR i_wbs_3_o_ack;
    o_wbm_1_i_ack       <= s_ack AND s_wbm_1_bg;
    o_wbm_2_i_ack       <= s_ack AND s_wbm_2_bg;
    -- rty
    s_rty <= i_wbs_1_o_rty OR i_wbs_2_o_rty OR i_wbs_3_o_rty;
    o_wbm_1_i_rty       <= s_rty AND s_wbm_1_bg;
    o_wbm_2_i_rty       <= s_rty AND s_wbm_2_bg;
    -- err
    s_err <= i_wbs_1_o_err OR i_wbs_2_o_err OR i_wbs_3_o_err;
    o_wbm_1_i_err       <= s_err AND s_wbm_1_bg;
    o_wbm_2_i_err       <= s_err AND s_wbm_2_bg;
  END BLOCK mux;

END ARCHITECTURE rtl;
